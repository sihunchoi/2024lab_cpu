// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define MEM_PATH mem
