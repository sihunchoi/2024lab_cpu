// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
//`define RF_PATH   CPU.icpu.i_datapath.rf
`define MEM_PATH mem
